// DO NOT SYNTHESIZE FILE
// This file is just a place holder for the IDE to detect the Vivado-generated IP core

module clk_wiz_golden_test (
    // Clock out ports
    output logic clk_out1,

    // Status and control signals
    input logic reset,
    output logic locked,

    // Clock in ports
    input logic clk_in1
);

endmodule
