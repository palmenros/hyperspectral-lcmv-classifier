// DO NOT SYNTHESIZE FILE
// This file is just a place holder for the IDE to detect the Vivado-generated IP core

module test_rom_w_1 (
    input logic clka,
    input logic[5:0] addra,
    output logic[31:0] douta
);

endmodule