// DO NOT SYNTHESIZE FILE
// This file is just a place holder for the IDE to detect the Vivado-generated IP core

module fp_adder_32_11 (
    input logic aclk,
    input logic aresetn,

    input logic s_axis_a_tvalid,
    input logic [31 : 0] s_axis_a_tdata,
    
    input logic s_axis_b_tvalid,
    input logic [31 : 0] s_axis_b_tdata,

    output logic m_axis_result_tvalid,
    output logic [31 : 0] m_axis_result_tdata
);
endmodule