// DO NOT SYNTHESIZE FILE
// This file is just a place holder for the IDE to detect the Vivado-generated IP core

module blk_mem_32_3 (
  input logic clka,
  input logic ena,
  input logic [0:0] wea,
  input logic [1:0] addra,
  input logic [31:0] dina,

  input logic clkb,
  input logic enb,
  input logic[1:0] addrb,
  output logic[31:0] doutb
);
endmodule