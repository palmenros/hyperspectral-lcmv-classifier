// DO NOT SYNTHESIZE FILE
// This file is just a place holder for the IDE to detect the Vivado-generated IP core

module uint32_to_float
(
  input logic aclk,
  input logic aresetn,
  input logic s_axis_a_tvalid,
  input logic[31:0] s_axis_a_tdata,
  output logic m_axis_result_tvalid,
  output logic[31:0] m_axis_result_tdata
);

endmodule